module Slave(input MOSI,);

endmodule
