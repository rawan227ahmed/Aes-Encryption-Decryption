module SPI();


endmodule
