module Inv_Mix_Columns(in,out);
input [0:127]in;
output [0:127]out;
/////////////////////////////////////////////////
function [0:7]multiply2;
input [0:7]x;
begin
if(x[0]==1)
multiply2=((x<<1)^8'h1b);
else
multiply2=x<<1;
end
endfunction 
////////////////////////////////////////////////
function [0:7]multiplye;  //e=8+4+1
input[0:7]x;
begin
multiplye=multiply2(multiply2(x))^multiply2(multiply2(multiply2(x)))^multiply2(x);
end
endfunction
/////////////////////////////////////////////////
function [0:7]multiplyd;   //d=8+2+1
input[0:7]x;
begin
multiplyd=multiply2(multiply2(x))^multiply2(multiply2(multiply2(x)))^x;
end
endfunction
//////////////////////////////////////////////////
function [0:7]multiplyb;   //
input[0:7]x;
begin
multiplyb=multiply2(multiply2(multiply2(x)))^multiply2(x)^x;
end
endfunction
//////////////////////////////////////////////////
function [0:7]multiply9;
input[0:7]x;
begin
multiply9=multiply2(multiply2(multiply2(x)))^x;
end
endfunction
//////////////////////////////////////////////////
genvar i;
generate
for(i=0;i<4;i=i+1)begin
assign out[(32*i)+:8]=multiplye(in[(32*i)+:8])^multiplyb(in[(32*i+8)+:8])^multiplyd(in[(32*i+16)+:8])^multiply9(in[(32*i+24)+:8]);
assign out[(32*i+8)+:8]=multiply9(in[(32*i)+:8])^multiplye(in[(32*i+8)+:8])^multiplyb(in[(32*i+16)+:8])^multiplyd(in[(32*i+24)+:8]);
assign out[(32*i+16)+:8]=multiplyd(in[(32*i)+:8])^multiply9(in[(32*i+8)+:8])^multiplye(in[(32*i+16)+:8])^multiplyb(in[(32*i+24)+:8]);
assign out[(32*i+24)+:8]=multiplyb(in[(32*i)+:8])^multiplyd(in[(32*i+8)+:8])^multiply9(in[(32*i+16)+:8])^multiplye(in[(32*i+24)+:8]);
end
endgenerate
endmodule 